
//package to define the scalable parameters
package p4_adder_pkg;

   parameter int nbit           = 32;
   parameter int nbit_per_block = 4;

endpackage
