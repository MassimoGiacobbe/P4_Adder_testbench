
//package to define the scalable parameters
package p4_pkg;

   parameter int nbit           = 32;
   parameter int nbit_per_block = 4;
   parameter int nTrans         = 5;
endpackage
